---------------------------------------------------------------------------------------------------
-- Copyright (c) 2025 Stefan Stähli
---------------------------------------------------------------------------------------------------

---------------------------------------------------------------------------------------------------
-- Description
---------------------------------------------------------------------------------------------------
-- This entity implements the Clark-PArke and D/Q transformed rquired for
-- field-oriented control (FOC).

---------------------------------------------------------------------------------------------------
-- Libraries
---------------------------------------------------------------------------------------------------
library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
  use IEEE.MATH_REAL.ALL;

library olo;
  use olo.en_cl_fix_pkg.all;
  use olo.olo_fix_pkg.all;

---------------------------------------------------------------------------------------------------
-- Entity Declaration
---------------------------------------------------------------------------------------------------
entity abc2dq is
    generic ( 
        DataWidth_g : natural
    );    
    port (
        -- Control Signals
        Clk         : in    std_logic;
        Rst         : in    std_logic;

        -- Modulator Inputs
        Sine        : in    std_logic_vector(DataWidth_g-1 downto 0);
        Cosine      : in    std_logic_vector(DataWidth_g-1 downto 0);
        -- ABC Inputs
        Strobe      : in    std_logic; -- new sample available
        A           : in    std_logic_vector(DataWidth_g-1 downto 0);
        B           : in    std_logic_vector(DataWidth_g-1 downto 0);
        C           : in    std_logic_vector(DataWidth_g-1 downto 0);
        -- DQ Outputs
        Valid       : out   std_logic; -- output data valid
        D           : out   std_logic_vector(DataWidth_g-1 downto 0);
        Q           : out   std_logic_vector(DataWidth_g-1 downto 0);
        DC          : out   std_logic_vector(DataWidth_g-1 downto 0)
    );
end abc2dq;

---------------------------------------------------------------------------------------------------
-- Architecture Declaration
---------------------------------------------------------------------------------------------------
architecture rtl of abc2dq is

    -- *** Constants ***
    constant FixFormat_c : FixFormat_t := (1, 0, DataWidth_g-1);
    constant FixFormatInt_c : FixFormat_t := cl_fix_add_fmt(FixFormat_c, FixFormat_c);
    
    constant cMtxPrescaler : real := 2.0/3.0; -- 2/3

    constant MtxCP11_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (           1.0), FixFormat_c); -- = 2/3
    constant MtxCP12_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (          -0.5), FixFormat_c); -- = -1/3
    constant MtxCP13_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (          -0.5), FixFormat_c); -- = -1/3
    constant MtxCP21_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (           0.0), FixFormat_c); -- = 0
    constant MtxCP22_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * ( sqrt(3.0)/2.0), FixFormat_c); -- = srt(3)/3
    constant MtxCP23_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (-sqrt(3.0)/2.0), FixFormat_c); -- = -sqrt(3)/3    
    constant MtxCP31_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (           0.5), FixFormat_c); -- = 1/3
    constant MtxCP32_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (           0.5), FixFormat_c); -- = 1/3
    constant MtxCP33_c : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0) := cl_fix_from_real(cMtxPrescaler * (           0.5), FixFormat_c); -- = 1/3

    constant NumStages_c : integer := 3; -- processing takes 3 pipeline stages (Valid on 4th edge after strobe)
    
    type SummandArray_t is array (0 to 2) of std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);

    type TwoProcess_r is record
        Sine : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        Cosine : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        Alpha : SummandArray_t;
        AlphaSum : std_logic_vector(cl_fix_width(FixFormatInt_c)-1 downto 0);
        Beta : SummandArray_t;
        BetaSum : std_logic_vector(cl_fix_width(FixFormatInt_c)-1 downto 0);
        Gamma : SummandArray_t;
        GammaSum : std_logic_vector(cl_fix_width(FixFormatInt_c)-1 downto 0);
        MtxDQ11 : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        MtxDQ12 : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        MtxDQ21 : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        MtxDQ22 : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        Valid : std_logic_vector(NumStages_c-1 downto 0);
        D : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        Q : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
        DC : std_logic_vector(cl_fix_width(FixFormat_c)-1 downto 0);
    end record;

    signal r, r_next : TwoProcess_r;

begin

    -----------------------------------------------------------------------------------------------
    -- Combinatorial Proccess
    -----------------------------------------------------------------------------------------------
    p_combinatorial: process(all) is
        variable v : TwoProcess_r;
    begin
        -- *** hold variables stable ***
        v := r;

        -- *** Default Values ***
        v.Sine := Sine;
        v.Cosine := Cosine;

        -- clarke transform (pipeline stage 1)
        v.Alpha(0) := cl_fix_mult(MtxCP11_c, FixFormat_c, A, FixFormat_c, FixFormat_c);
        v.Alpha(1) := cl_fix_mult(MtxCP12_c, FixFormat_c, B, FixFormat_c, FixFormat_c);
        v.Alpha(2) := cl_fix_mult(MtxCP13_c, FixFormat_c, C, FixFormat_c, FixFormat_c);

        v.Beta(0)  := cl_fix_mult(MtxCP21_c, FixFormat_c, A, FixFormat_c, FixFormat_c);
        v.Beta(1)  := cl_fix_mult(MtxCP22_c, FixFormat_c, B, FixFormat_c, FixFormat_c);
        v.Beta(2)  := cl_fix_mult(MtxCP23_c, FixFormat_c, C, FixFormat_c, FixFormat_c);
        
        v.Gamma(0) := cl_fix_mult(MtxCP31_c, FixFormat_c, A, FixFormat_c, FixFormat_c);
        v.Gamma(1) := cl_fix_mult(MtxCP32_c, FixFormat_c, B, FixFormat_c, FixFormat_c);
        v.Gamma(2) := cl_fix_mult(MtxCP33_c, FixFormat_c, C, FixFormat_c, FixFormat_c);

        -- simplified park transform (pipeline stage 2)
        v.MtxDQ11 := cl_fix_resize(r.Cosine, FixFormat_c, FixFormat_c);
        v.MtxDQ12 := cl_fix_resize(r.Sine, FixFormat_c, FixFormat_c);
        v.MtxDQ21 := cl_fix_neg(r.Sine, FixFormat_c, FixFormat_c, saturate => Sat_s);
        v.MtxDQ22 := cl_fix_resize(r.Cosine, FixFormat_c, FixFormat_c);

        -- clarke transform sumup (pipeline stage 2)
        v.AlphaSum := cl_fix_add(
            cl_fix_add(
                r.Alpha(0), FixFormat_c,
                r.Alpha(1), FixFormat_c,
                FixFormatInt_c), FixFormatInt_c,
            r.Alpha(2), FixFormat_c,
            FixFormatInt_c);
            
        v.BetaSum  := cl_fix_add(
            cl_fix_add(
                r.Beta(0), FixFormat_c,
                r.Beta(1), FixFormat_c,
                FixFormatInt_c), FixFormatInt_c,
            r.Beta(2), FixFormat_c,
            FixFormatInt_c);

        v.GammaSum := cl_fix_add(
            cl_fix_add(
                r.Gamma(0), FixFormat_c,
                r.Gamma(1), FixFormat_c,
                FixFormatInt_c), FixFormatInt_c,
            r.Gamma(2), FixFormatInt_c,
            FixFormatInt_c);

        -- calc outputs (pipeline stage 3)
        v.D := cl_fix_add(
            cl_fix_mult(r.MtxDQ11, FixFormat_c, r.AlphaSum, FixFormatInt_c, FixFormatInt_c), FixFormatInt_c, 
            cl_fix_mult(r.MtxDQ12, FixFormat_c, r.BetaSum, FixFormatInt_c, FixFormatInt_c), FixFormatInt_c,
            FixFormat_c, saturate => Sat_s);
        v.Q := cl_fix_add(
            cl_fix_mult(r.MtxDQ21, FixFormatInt_c, r.AlphaSum, FixFormatInt_c, FixFormatInt_c), FixFormatInt_c, 
            cl_fix_mult(r.MtxDQ22, FixFormatInt_c, r.BetaSum, FixFormatInt_c, FixFormatInt_c), FixFormatInt_c, 
            FixFormat_c, saturate => Sat_s);
        v.DC := cl_fix_resize(
            r.GammaSum, FixFormatInt_c,
            FixFormat_c, saturate => Sat_s
        );

        v.Valid := r.Valid(r.Valid'left-1 downto 0) & Strobe;

        r_next <= v;
    end process p_combinatorial;

    -----------------------------------------------------------------------------------------------
    -- Outputs
    -----------------------------------------------------------------------------------------------
    Valid <= r.Valid(r.Valid'left);
    D <= r.D;
    Q <= r.Q;
    DC <= r.DC;

    -----------------------------------------------------------------------------------------------
    -- Sequential Proccess
    -----------------------------------------------------------------------------------------------
    p_seq : process (Clk) is
    begin
        if rising_edge(Clk) then
            r <= r_next;
            if Rst = '1' then
                r.Valid <= (others => '0');
                r.D <= (others => '0');
                r.Q <= (others => '0');
                r.DC <= (others => '0');
            end if;
        end if;
    end process;

end architecture;